
// Behavioural models for supply filter capacitors

module FilterCapCellDig (
        inout VDD,
        inout GND);
endmodule

module FilterCapDig_2x2 (
        inout VDD,
        inout GND);
endmodule

module FilterCap_DVDD_1 (
        inout VDD,
        inout GND);
endmodule

module FilterCap_DVDD_2 (
        inout VDD,
        inout GND);
endmodule

module FilterCap_DVDD_3 (
        inout VDD,
        inout GND);
endmodule


