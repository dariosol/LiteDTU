module IO_CORNER (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);
endmodule

