module IO_FILLER20 (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);

endmodule

module IO_FILLER10 (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);

endmodule

module IO_FILLER5 (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);

endmodule

module IO_FILLER1 (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);

endmodule

module IO_FILLER05 (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);

endmodule

module IO_FILLER0005 (
	inout VDD,
	inout VSS,
	inout VDDPST,
	inout VSSPST);

endmodule

